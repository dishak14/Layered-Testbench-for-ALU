interface intf();
  logic [7:0] a;
  logic[7:0] b;
  logic [1:0] s;
  logic [8  :0] y;
endinterface
